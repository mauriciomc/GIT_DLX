library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity INS_MEM is
	generic (N : integer);
	port (RST : in std_logic;
			CLK : in std_logic;
			address : in std_logic_vector (6 downto 0);
			data : out std_logic_vector (N-1 downto 0));
		
end INS_MEM;

architecture Structural of INS_MEM is
type Rom_Array is array (0 to 127) of std_logic_vector(7 downto 0);
signal content : Rom_Array;

begin

MEM: process (address)
	variable index : integer := 0;
	begin		
		
		Content <= ("00100000","00000001","00000000","00100000",  --0  addi $1  $0  32    
						"00100000","00010100","00000000","10001101",  --4  addi $20 $0  141
						"00000000","00110100","00101000","00100000",  --8  add  $5  $20  $1
						"10101100","00000001","00000000","00000101",  --12  sw  $1  MEM[5]
						"00001000","00000000","00000000","00001110",  --16 jmp  14*4 = 56
						"00100000","00000000","00000000","00000000",  --20 nop		 
						"00100000","00000000","00000000","00000000",  --24 nop		 
						"00100000","00000000","00000000","00000000",  --28 nop	
						"00100000","00000000","00000000","00000000",  --32 nop		 
						"00000011","11111111","11111000","00001000",  --36 jr  $31 
						"00100000","00000000","00000000","00000000",  --40 nop		 
						"00100000","00000000","00000000","00000000",  --44 nop		 
						"00100000","00000000","00000000","00000000",  --48 nop	
						"00100000","00000000","00000000","00000000",  --52 nop		 
						"10001100","00001000","00000000","00000101",  --56  lw  $8  MEM[5]
						"00000000","00100001","11000000","00011000",  --60  mul $24 $1  $1
						"00100000","00111101","00000000","01000000",  --64 addi $29 $1  64 
						"00100000","00000000","00000000","00000000",  --68 nop		 
						"00100000","00000000","00000000","00000000",  --72 nop		 
						"00100000","00000000","00000000","00000000",  --76 nop		 
						"00100000","00000000","00000000","00000000",  --80 nop		 
						"00001100","00000000","00000000","00001001",  --84 jal 36 = 9*4
   					"00100000","00000000","00000000","00000000",  --88 nop		 
						"00100000","00000000","00000000","00000000",  --92 nop		 
						"00100000","00000000","00000000","00000000",  --96 nop		 
						"00100000","00000000","00000000","00000000",  --100 nop		 
						"00000000","00011101","11101001","10000011",  --104 sra  $29 6
						"00000000","00101000","01000000","00011000",  --108 mul  $8 $8 $1 
						"00010100","00000101","11111111","11110000",  --112 bne  $5 -4 (= NPC-8)
						"00100000","00000000","00000000","00000000",  --116 nop		 
						"00100000","00000000","00000000","00000000",  --120 nop		 
						"00100000","00000000","00000000","00000000"); --124 nop		 
				
				
		index := conv_integer(unsigned(address));
		data <= content(index) & content(index+1) & content(index+2) & content(index+3);

	end process;
end Structural;

-- Some testable programs -- Without Hazard RAW control

--					  ("00100000","00000001","00000000","00000101", --0  addi $1 $0 5
--						"00100000","00000000","00000000","00000000", --4  nop
--						"00100000","00000000","00000000","00000000", --8  nop
--						"00100000","00000000","00000000","00000000", --12 nop
--						"00100000","00000000","00000000","00000000", --16 nop
--						"00011100","00100000","00000000","00010000", --20 bgtz $1 16(+NPC=40)
--						"00100000","00100001","11111111","11111111", --24 addi $1 $1 -1
--						"00100000","00000000","00000000","00000000", --28 nop
--						"00100000","00000000","00000000","00000000", --32 nop
--						"00100000","00000000","00000000","00000000", --36 nop
--						"00100000","00000000","00000000","00000000", --40 nop
--						"10101100","00100000","00000000","00000100", --44 sw $1 4
--						"00010100","00100000","11111111","11110010", --48 bne $1 -28(+NPC=24)
--		            "00001000","00000000","00000000","00000000");--52 jmp 0


--PC=0           
		-- addi 			   "001000"   To perform a move to register 
		-- (Rs unuse		"00000")
		-- in R[1] (value: 0)"00001"
		-- the immediate 5  "0000000000000101"
		
--PC=4
		-- addi 				     "001000"   To perform a NOP
		-- (Rs unused			  "00000" )
		-- in R[0]  (value: 0) "00000"
		-- the immediate 0	  "0000000000000000" 

--PC=8
		-- addi 				     "001000"   To perform a NOP
		-- (Rs unused			  "00000" )
		-- in R[0]  (value: 0) "00000"
		-- the immediate 0	  "0000000000000000" 

--PC=12
		-- addi 				     "001000"   To perform a NOP
		-- (Rs unused			  "00000" )
		-- in R[0]  (value: 0) "00000"
		-- the immediate 0	  "0000000000000000" 

--PC=16
		-- addi 				     "001000"   To perform a NOP
		-- (Rs unused			  "00000" )
		-- in R[0]  (value: 0) "00000"
		-- the immediate 0	  "0000000000000000" 

--PC=20
		-- bgtz 				     "000111"   Branch if greater than zero
		-- (Rs unused			  "00001")
		-- in R[0]  (value: 0) "00000"
		-- the immediate 28	  "0000000000011100" 

--PC=24
		-- addi 				     "001000"   To perform a NOP
		-- (Rs unused			  "00001" )
		-- in R[0]  (value: 0) "00001"
		-- the immediate -1	  "1111111111111110" 

--PC=28
		-- addi 				     "001000"   To perform a NOP
		-- (Rs unused			  "00000" )
		-- in R[0]  (value: 0) "00000"
		-- the immediate 0	  "0000000000000000" 

--PC=32
		-- addi 				     "001000"   To perform a NOP
		-- (Rs unused			  "00000" )
		-- in R[0]  (value: 0) "00000"
		-- the immediate 0	  "0000000000000000" 

--PC=36
		-- addi 				     "001000"   To perform a NOP
		-- (Rs unused			  "00000" )
		-- in R[0]  (value: 0) "00000"
		-- the immediate 0	  "0000000000000000" 

--PC=40
		-- addi 				     "001000"   To perform a NOP
		-- (Rs unused			  "00000" )
		-- in R[0]  (value: 0) "00000"
		-- the immediate 0	  "0000000000000000" 

--PC=44
		-- sw 				     "101011"   Store word
		-- (Rs unused			  "00000" )
		-- in R[1]             "00001"
		-- the immediate 20    "0000000000010100" 

--PC=48
		-- bne 				     "000101"   Branch if Rs != 0
		-- (Rs unused			  "00001" )
		-- in R[0]  (value: 0) "00000"
		-- the immediate 0	  "0000000000011000" 
--PC=52
		-- jmp 				     "000010"   To perform a NOP
		-- target 0       	  "0000000000000000" 

